interface dff_if(input logic clk);
    logic rst_n;
    logic d;
    logic q;
endinterface